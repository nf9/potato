// Verilog netlist created by TD v4.5.12562
// Tue Jul 30 23:36:08 2019

`timescale 1ns / 1ps
module instruction_rom  // al_ip/bram.v(14)
  (
  addra,
  clka,
  rsta,
  doa
  );

  input [10:0] addra;  // al_ip/bram.v(18)
  input clka;  // al_ip/bram.v(19)
  input rsta;  // al_ip/bram.v(20)
  output [31:0] doa;  // al_ip/bram.v(16)


  assign doa[31] = doa[3];
  assign doa[30] = doa[2];
  assign doa[29] = doa[1];
  assign doa[28] = doa[0];
  assign doa[27] = doa[3];
  assign doa[26] = doa[2];
  assign doa[25] = doa[1];
  assign doa[24] = doa[0];
  assign doa[23] = doa[3];
  assign doa[22] = doa[2];
  assign doa[21] = doa[1];
  assign doa[20] = doa[0];
  assign doa[19] = doa[3];
  assign doa[18] = doa[2];
  assign doa[17] = doa[1];
  assign doa[16] = doa[0];
  assign doa[15] = doa[3];
  assign doa[14] = doa[2];
  assign doa[13] = doa[1];
  assign doa[12] = doa[0];
  assign doa[11] = doa[3];
  assign doa[10] = doa[2];
  assign doa[9] = doa[1];
  assign doa[8] = doa[0];
  assign doa[7] = doa[3];
  assign doa[6] = doa[2];
  assign doa[5] = doa[1];
  assign doa[4] = doa[0];
  EG_PHY_CONFIG #(
    .DONE_PERSISTN("ENABLE"),
    .INIT_PERSISTN("ENABLE"),
    .JTAG_PERSISTN("DISABLE"),
    .PROGRAMN_PERSISTN("DISABLE"))
    config_inst ();
  // address_offset=0;data_offset=0;depth=2048;width=4;num_section=1;width_per_section=4;section_size=32;working_depth=2048;working_width=4;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("4"),
    .DATA_WIDTH_B("4"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_2048x32_sub_000000_000 (
    .addra({addra,2'b11}),
    .clka(clka),
    .dia({open_n69,open_n70,open_n71,open_n72,open_n73,4'b0000}),
    .rsta(rsta),
    .doa({open_n88,open_n89,open_n90,open_n91,open_n92,doa[3:0]}));

endmodule 

